shared/keyscans.vh